module counter_tb;
  
  bit clk, reset_n, up_down;
  bit 
  
endmodule
